/*
Header file containing all decodings of the command hex encoding
*/

`define UPDATE_SCORE_COMMAND 8'b0001xxxx
`define CHANGE_SCREEN_COMMAND 8'b0010xxxx // We might not actually need this
`define COLOR_COMMAND 8'b1000xxxx
