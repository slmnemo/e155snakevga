/*
Module to decode SPI commands
*/

module command_decoder (
    
);