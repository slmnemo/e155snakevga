/*
Define file for VGA timings, fetch timings, and 


*/
`define RISETIMECORRECTION 0

`define HACTIVE 640
`define HFRONTPORCH 16
`define HSYNCPULSE 96
`define HBACKPORCH 48
`define HFULLSCAN (`HACTIVE+`HFRONTPORCH+`HSYNCPULSE+`HBACKPORCH)

`define VACTIVE 480
`define VFRONTPORCH 11
`define VSYNCPULSE 2
`define VBACKPORCH 32
`define VFULLSCAN (`VACTIVE+`VFRONTPORCH+`VSYNCPULSE+`VBACKPORCH)

`define HFETCHNEXTLINE 20
`define HFETCH `HFULLSCAN - `HFETCHNEXTLINE - 1

// Offsets for number positions

`define ONES_X_OFFSET 639
`define TENS_X_OFFSET 619
`define HUNS_X_OFFSET 599

`define ONES_Y_OFFSET 479
`define TENS_Y_OFFSET 479
`define HUNS_Y_OFFSET 479


