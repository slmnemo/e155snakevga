/*
Header file containing all decodings of the command hex encoding
*/

`define UPDATE_SCORE_COMMAND 8'b0001????
`define CHANGE_SCREEN_COMMAND 8'b0010???? // We might not actually need this
`define COLOR_COMMAND 8'b1000????
